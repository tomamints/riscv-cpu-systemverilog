import eei::*;
import corectrl::*;

module csrunit (
	input  logic clk,
	input  logic rst,
	input  logic valid,
	input  Addr  pc,
	input  Inst  inst_bits,
	input  InstCtrl ctrl,
	input  ExceptionInfo expt_info,
	input  logic [4:0]  rd_addr,
	input  logic [11:0] csr_addr,
	input  logic [4:0]  rs1_addr,
	input  UIntX rs1_data,
	input  logic can_intr,
	output UIntX rdata,
	output PrivMode mode,
	output logic raise_trap,
	output Addr  trap_vector,
	output logic trap_return,
	input  UInt64  minstret,
	aclint_if.slave aclint
);

//WMASK determines which bit can change or not. WARL can write anything but read legal.
	localparam UIntX MSTATUS_WMASK = UIntX'('h0000_0000_0060_19aa) ;
	localparam UIntX MTVEC_WMASK  = 'hffff_ffff_ffff_fffd; //MTVECは[1:0]はMODE設定
	localparam UIntX MEDELEG_WMASK  = 'hffff_ffff_ffff_f7ff;
	localparam UIntX MIDELEG_WMASK  = UIntX'('h0000_0000_0000_0222);
	localparam UIntX MCOUNTEREN_WMASK  = UIntX'('h0000_0000_0000_0007);
	localparam UIntX MSCRATCH_WMASK = 'hffff_ffff_ffff_ffff;
	localparam UIntX MEPC_WMASK   = 'hffff_ffff_ffff_fffe;
	localparam UIntX MCAUSE_WMASK = 'hffff_ffff_ffff_ffff;
	localparam UIntX MTVAL_WMASK  = 'hffff_ffff_ffff_ffff;
	localparam UIntX MIP_WMASK  = UIntX'('h0000_0000_0000_0222);
	localparam UIntX MIE_WMASK  = UIntX'('h0000_0000_0000_02aa);

	localparam UIntX SSTATUS_WMASK  = UIntX'('h0000_0000_0000_0122);
	localparam UIntX SIE_WMASK      = UIntX'('h0000_0000_0000_0222);
	localparam UIntX SCOUNTEREN_WMASK  = UIntX'('h0000_0000_0000_0007);
	localparam UIntX STVEC_WMASK  = 'hffff_ffff_ffff_fffd;
	localparam UIntX SSCRATCH_WMASK = 'hffff_ffff_ffff_ffff;
	localparam UIntX SEPC_WMASK   = 'hffff_ffff_ffff_fffe;
	localparam UIntX SCAUSE_WMASK = 'hffff_ffff_ffff_ffff;
	localparam UIntX STVAL_WMASK  = 'hffff_ffff_ffff_ffff;


	//read masks
	localparam UIntX SSTATUS_RMASK  = UIntX'('h8000_0003_018f_e762);


	//CSRR(W|S|C)かどうか
	logic is_wsc;
	assign is_wsc = ctrl.is_csr && ctrl.funct3[1:0] != 0;

	logic is_mret;
	assign is_mret = (inst_bits == 32'h30200073);

	logic is_sret;
	assign is_sret = (inst_bits == 32'h10200073);

	logic is_wfi;
	assign is_wfi = (inst_bits == 32'h10500073);

	// will_not_write_csr: CSRRSI / CSRRCI で rs1=0 のとき → 読み取り専用動作
	logic will_not_write_csr;
	assign will_not_write_csr =
		((ctrl.funct3[1:0] == 2'b10) || (ctrl.funct3[1:0] == 2'b11))
		&& (rs1_addr == 5'd0);

	// expt_write_readonly_csr: 書き込み系で、書き込み禁止CSRにアクセスしたとき
	logic expt_write_readonly_csr;
	assign expt_write_readonly_csr =
		(is_wsc && !will_not_write_csr && (csr_addr[11:10] == 2'b11));

	logic expt_csr_priv_violation;
	assign expt_csr_priv_violation = is_wsc && (csr_addr[9:8] > mode);

	logic expt_zicntr_priv;
	logic zicntr_denied_S;
	assign zicntr_denied_S =
		(csr_addr == CYCLE)   ? !mcounteren[0] :
		(csr_addr == TIME)    ? !mcounteren[1] :
		(csr_addr == INSTRET) ? !mcounteren[2] :
										1'b0;

	logic zicntr_denied_U =
		(csr_addr == CYCLE)   ? !scounteren[0] :
		(csr_addr == TIME)    ? !scounteren[1] :
		(csr_addr == INSTRET) ? !scounteren[2] :
										1'b0;

	assign expt_zicntr_priv =
		is_wsc &&
		(mode <= S &&
		zicntr_denied_S ||
		zicntr_denied_U);

	logic expt_trap_return_priv;
	assign expt_trap_return_priv = (is_mret && mode < M) || (is_sret && mode < S || (mode == S && mstatus_tsr));
	//attempt to execute trap return instruction in low privilege level

	//CSR register create
	UIntX misa;
	assign misa = {
    2'd2,                                         // MISAの最上位2ビット (MISA[XLEN-1:XLEN-2])
    1'b0,                                         // 次の1ビット
    {(XLEN - 2 - 1 - 26){1'b0}},                  // 'repeat XLEN - 28' に相当する0ビットの繰り返し
                                                  // (XLEN - 28) = XLEN - (2 + 1 + 25) ではなく、
                                                  // XLEN - (2 + 1 + 26) = XLEN - 29 が正しいため、
                                                  // XLEN - 2 - 1 - 26 = XLEN - 29 で計算します。
    26'b00000101000001000100000101                // MISAの最下位26ビット
	};

	UIntX mhartid = 0;
	UIntX mstatus, mtvec, mideleg, mie, mip, mip_reg, mscratch, mepc, mcause, mtval;
	UInt32 mcounteren;
	UInt64 mcycle, medeleg;

	assign mip = mip_reg | {
		{(XLEN - 12){1'b0}},
		1'b0, // MEIP
		1'b0, // 0
		1'b0, // SEIP
		1'b0, // 0
		aclint.mtip, // MTIP
		1'b0, // 0
		1'b0, // STIP
		1'b0, // 0
		aclint.msip, //MSIP
		1'b0, // 0
		1'b0, // SSIP
		1'b0 // 0
	};



	//mstatus bits

	logic mstatus_tsr;
	assign mstatus_tsr = mstatus[22];

	PrivMode mstatus_mpp;
	assign mstatus_mpp = PrivMode'(mstatus[12:11]);

	PrivMode mstatus_spp;
	assign mstatus_spp = (mstatus[8]) ? S : U;

	logic mstatus_mpie;
	assign mstatus_mpie = mstatus[7];

	logic mstatus_mie;
	assign mstatus_mie = mstatus[3];

	logic mstatus_sie;
	assign mstatus_sie = mstatus[1];

	//Supevisor mode CSR
	UIntX  sstatus , stvec, sscratch, sip, sie, sepc, scause, stval;
	assign sstatus = mstatus & SSTATUS_RMASK;
	UInt32 scounteren;

	assign sip = mip & mideleg;

	//Interrupt to M-mode
	UIntX interrupt_pending_mmode;
	assign interrupt_pending_mmode = mip & mie & ~mideleg;
	logic raise_interrupt_mmode;
	assign raise_interrupt_mmode = (mode != M || mstatus_mie) && interrupt_pending_mmode != 0;

	UIntX interrupt_cause_mmode;
	assign interrupt_cause_mmode =
		interrupt_pending_mmode[3] ? MACHINE_SOFTWARE_INTERRUPT :
		interrupt_pending_mmode[7] ? MACHINE_TIMER_INTERRUPT :
		interrupt_pending_mmode[9] ? SUPERVISOR_EXTERNAL_INTERRUPT :
		interrupt_pending_mmode[1] ? SUPERVISOR_SOFTWARE_INTERRUPT :
		interrupt_pending_mmode[5] ? SUPERVISOR_TIMER_INTERRUPT :
							UIntX'(0);

	//Interrupt to S-mode
	UIntX interrupt_pending_smode;
	assign interrupt_pending_smode = sip & sie;
	logic raise_interrupt_smode;
	assign raise_interrupt_smode = (mode < S || (mode == S && mstatus_sie)) && interrupt_pending_smode != 0;

	UIntX interrupt_cause_smode;
	assign interrupt_cause_smode =
		interrupt_pending_smode[9] ? SUPERVISOR_EXTERNAL_INTERRUPT :
		interrupt_pending_smode[1] ? SUPERVISOR_SOFTWARE_INTERRUPT :
		interrupt_pending_smode[5] ? SUPERVISOR_TIMER_INTERRUPT :
							UIntX'(0);


		//Interrupt
	logic raise_interrupt;
	assign raise_interrupt = valid && can_intr && (raise_interrupt_mmode || raise_interrupt_smode);

	UIntX interrupt_cause;
	assign interrupt_cause = (raise_interrupt_mmode) ? interrupt_cause_mmode : interrupt_cause_smode;

	Addr interrupt_xtvec;
	assign interrupt_xtvec = (interrupt_mode == M) ? mtvec: stvec;

	Addr interrupt_vector;
	assign interrupt_vector = (interrupt_xtvec[0] == 0) ? {interrupt_xtvec[XLEN-1 : 2], 2'b0} : { (interrupt_xtvec[XLEN-1:2] + interrupt_cause[XLEN-1-2:0]),2'b0}; //vectored

	PrivMode interrupt_mode;
	assign interrupt_mode = (raise_interrupt_mmode) ? M : S ;

	//Exception
	logic raise_expt;
	assign raise_expt = valid && (expt_info.valid || expt_write_readonly_csr || expt_csr_priv_violation || expt_zicntr_priv || expt_trap_return_priv);
	UIntX expt_cause ;
	always_comb begin
		if(expt_info.valid) begin
			expt_cause = expt_info.cause;
		end else if (expt_write_readonly_csr) begin
			expt_cause = ILLEGAL_INSTRUCTION;
		end else if (expt_csr_priv_violation) begin
			expt_cause = ILLEGAL_INSTRUCTION;
		end else if (expt_zicntr_priv) begin
			expt_cause = ILLEGAL_INSTRUCTION;
		end else if (expt_trap_return_priv) begin
			expt_cause = ILLEGAL_INSTRUCTION;
		end else begin
			expt_cause = '0;
		end
	end

	UIntX expt_value;
	always_comb begin
		if (expt_info.valid)begin
			expt_value = expt_info.value;
		end else if (expt_cause == ILLEGAL_INSTRUCTION) begin
			expt_value = { {(XLEN - $bits(Inst)){1'b0}}, inst_bits };
		end else begin
			expt_value = '0;
		end
	end

	Addr expt_xtvec;
	assign expt_xtvec = (expt_mode == M) ? mtvec : stvec;

	Addr expt_vector;
	assign expt_vector = {expt_xtvec[XLEN-1 : 2], 2'b0};

	PrivMode expt_mode;
	assign expt_mode = (mode == M || !medeleg[expt_cause[5:0]]) ? M : S;

	// Trap Return
	assign trap_return = valid && (is_mret || is_sret) && !raise_expt && !raise_interrupt;
	PrivMode trap_return_mode;
	assign trap_return_mode = (is_mret) ? mstatus_mpp : mstatus_spp;
	Addr trap_return_vector ;
	assign trap_return_vector = (is_mret) ? mepc : sepc;


	//Trap
	assign raise_trap  = raise_expt || raise_interrupt || trap_return;

	UIntX  trap_cause ;
	assign trap_cause =
    raise_expt      ? expt_cause :
    raise_interrupt ? interrupt_cause :
                      UIntX'(0);

	assign trap_vector =
		raise_expt      ? expt_vector :
		raise_interrupt ? interrupt_vector :
		trap_return     ? trap_return_vector :
						UIntX'(0);

	PrivMode trap_mode_next;
	assign trap_mode_next =
		raise_expt      ? expt_mode :
		raise_interrupt ? interrupt_mode :
		trap_return     ? trap_return_mode :
						  U;   // enum名は環境に合わせて



	UIntX wdata;
	UIntX wmask;

	logic [XLEN-1:0] wsource; //always_comb の外で定義

	always_comb begin
		// read
		case (csr_addr)
			MISA    : rdata = misa;
			MIMPID  : rdata = MACHINE_IMPLEMENTATION_ID;
			MHARTID : rdata = mhartid;
			MSTATUS : rdata = mstatus;
			MTVEC   : rdata = mtvec;
			MEDELEG   : rdata = medeleg;
			MIDELEG   : rdata = mideleg;
			MIP   : rdata = mip;
			MIE   : rdata = mie;
			MCOUNTEREN   : rdata = {{(XLEN-32){1'b0}},mcounteren};
			MCYCLE  : rdata = mcycle;
			MINSTRET: rdata = minstret;
			MSCRATCH: rdata = mscratch;
			MEPC    : rdata = mepc;
			MCAUSE  : rdata = mcause;
			MTVAL   : rdata = mtval;
			SSTATUS   : rdata = sstatus;
			SCOUNTEREN : rdata = {{(XLEN - 32){1'b0}}, scounteren};
			STVEC   : rdata = stvec;
			SEPC    : rdata = sepc;
			SCAUSE  : rdata = scause;
			STVAL   : rdata = stval;
			SIP     : rdata = sip;
			SIE     : rdata = sie & mideleg;
			CYCLE   : rdata = mcycle;
			TIME    : rdata = aclint.mtime;
			INSTRET : rdata = minstret;
			default       : rdata = 'x;
		endcase

		// write mask
		case (csr_addr)
			MSTATUS  : wmask = MSTATUS_WMASK;
			MTVEC    : wmask = MTVEC_WMASK;
			MEDELEG    : wmask = MEDELEG_WMASK;
			MIDELEG    : wmask = MIDELEG_WMASK;
			MIP      : wmask = MIP_WMASK;
			MIE      : wmask = MIE_WMASK;
			MCOUNTEREN : wmask = MCOUNTEREN_WMASK;
			MSCRATCH : wmask = MSCRATCH_WMASK;
			MEPC     : wmask = MEPC_WMASK;
			MCAUSE   : wmask = MCAUSE_WMASK;
			MTVAL    : wmask = MTVAL_WMASK;
			SSTATUS  : wmask = SSTATUS_WMASK;
			SCOUNTEREN : wmask = SCOUNTEREN_WMASK;
			STVEC : wmask = STVEC_WMASK;
			SSCRATCH : wmask = SSCRATCH_WMASK;
			SCAUSE : wmask = SCAUSE_WMASK;
			STVAL : wmask = STVAL_WMASK;
			SIE : wmask = SIE_WMASK & mideleg;
			default       : wmask = '0;
		endcase

		// wsource
		// (funct3[2] == 1 : immediate → rs1_addr is used)
		if (ctrl.funct3[2]) begin
			wsource = {{(XLEN-5){1'b0}}, rs1_addr};
		end else begin
			wsource = rs1_data;
		end

		// wdata (CSRRS, CSRRC, etc.)
		case (ctrl.funct3[1:0])
			2'b01:  wdata = wsource;            // CSRRW / CSRRWI
			2'b10:  wdata = rdata | wsource;    // CSRRS / CSRRSI
			2'b11:  wdata = rdata & ~wsource;   // CSRRC / CSRRCI
			default: wdata = 'x;
		endcase

		// apply write mask
		wdata = (wdata & wmask) | (rdata & ~wmask);
	end

	UIntX setssip;
	assign setssip = {{(XLEN - 2){1'b0}}, aclint.setssip, 1'b0 };

	Addr xepc;

	always_ff @(posedge clk or negedge rst) begin
		if (!rst) begin
			mode     <=  M;
			mstatus  <=  MSTATUS_UXL | MSTATUS_SXL;
			mtvec    <= '0;
			medeleg    <= '0;
			mideleg    <= '0;
			mie      <= '0;
			mip_reg  <= '0;
			mcounteren <= '0;
			mscratch <= '0;
			mcycle   <= '0;
			mepc     <= '0;
			mcause   <= '0;
			mtval    <= '0;
			scounteren <= '0;
			stvec <= '0;
			sscratch <= '0;
			sepc <= '0;
			scause <= '0;
			stval <= '0;
			sie <= '0;
		end else begin
			mcycle += 1;
			mip_reg |= setssip;
			if (valid) begin
				if (raise_trap) begin
					if (raise_expt || raise_interrupt) begin
						if (raise_expt)begin
							xepc = pc; //exception
						end else if (raise_interrupt && is_wfi) begin
							xepc = pc + 4;
						end else begin
							xepc = pc;
						end
						if (trap_mode_next == M) begin
							mepc <= xepc;
							mcause <= trap_cause;
							if (raise_expt) begin
								mtval <= expt_value;
							end
							//save mstatus.mie to mstatus.mpie
							//and set mstatus.mie = 0
							mstatus[7] <= mstatus[3];
							mstatus[3] <= 0;
							//save current priviledge level to mstatus.mpp
							mstatus[12:11] <= mode;
						end else begin
							sepc <= xepc;
							scause <= trap_cause;
							if (raise_expt) begin
								stval <= expt_value;
							end
							//save sstatus.sie to sstatus.spie
							//and set sstatus.sie = 0
							mstatus[5] <= mstatus[1];
							mstatus[1] <= 0;
							//save current privilege mode (S or U) to sstatus.spp
							mstatus[8] <= mode[0];
						end
					end else if (trap_return) begin
						if (is_mret) begin
							//save mstatus.mie to mstatus.mipe
							// and set mstatus.mie = 0
							mstatus[3] <= mstatus[7];
							mstatus[7] <= 0;
							// set mstatus.mpp = U (least priviledge level)
							mstatus[12:11] <= U;
						end else if (is_sret) begin
							//set sstatus.sie = sstatus.spie
							//    sstatus.spie = 0
							mstatus[1] <= mstatus[5];
							mstatus[5] <= 0;
							//set sstatus.spp <= U
							mstatus[8] <= 0;
						end
					end
					mode <= trap_mode_next;
				end else begin
					if (is_wsc) begin
						case (csr_addr) //これらはそれぞれのCSRレジスタにwdataを入れている。
							MSTATUS  : mstatus  <= validate_mstatus(mstatus, wdata);
							MTVEC    : mtvec    <= wdata;
							MEDELEG    : medeleg    <= wdata;
							MIDELEG   : mideleg    <= wdata;
							MIP      : mip_reg    <= (wdata & MIP_WMASK) | setssip;
							MIE      : mie      <= wdata & MIE_WMASK;
							MCOUNTEREN : mcounteren <= wdata[31:0];
							MSCRATCH : mscratch <= wdata;
							MEPC     : mepc     <= wdata;
							MCAUSE   : mcause   <= wdata;
							MTVAL    : mtval    <= wdata;
							SSTATUS  : mstatus  <= validate_mstatus(mstatus, wdata | mstatus & ~SSTATUS_WMASK);
							SCOUNTEREN : scounteren <= wdata[31:0];
							STVEC : stvec <= wdata;
							SSCRATCH : sscratch <= wdata;
							SEPC : sepc <= wdata;
							SCAUSE : scause <= wdata;
							STVAL : stval <= wdata;
							SIE : sie <= wdata;
							default  : /* do nothing */ ;
						endcase
					end
				end
			end
		end
	end
	function automatic UIntX validate_mstatus(
		input UIntX mstatus,
		input UIntX wdata
	);
		UIntX result;
		result = wdata;

		// MPP: only M(11) or U(00) allowed
		if (wdata[12:11] == 2'b10)
		begin
			result[12:11] = mstatus[12:11];
		end

		return result;
	endfunction
endmodule : csrunit
