import eei::*;

module dma_regs (
    input logic mmio_valid,
    input logic mmio_we,
);


endmodule
